LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY EECE381_NUMERIC_HEX IS
	PORT(
	   	NUM	: IN  STD_LOGIC_VECTOR(3 DOWNTO 0);	-- Number to be displayed
	   	SEG7	: OUT STD_LOGIC_VECTOR(6 DOWNTO 0)	-- Seven segment display to use
	);
END;


ARCHITECTURE BEHAVIOURAL OF EECE381_NUMERIC_HEX IS

	

BEGIN

	PROCESS (NUM)
	BEGIN
		CASE NUM IS
		WHEN "0000" => SEG7 <= "1000000";	-- 0
		WHEN "0001" => SEG7 <= "1111001";	-- 1
		WHEN "0010" => SEG7 <= "0100100";	-- 2
		WHEN "0011" => SEG7 <= "0110000";	-- 3
		WHEN "0100" => SEG7 <= "0011001";	-- 4
		WHEN "0101" => SEG7 <= "0010010";	-- 5
		WHEN "0110" => SEG7 <= "0000010";	-- 6
		WHEN "0111" => SEG7 <= "1111000";	-- 7
		WHEN "1000" => SEG7 <= "0000000";	-- 8
		WHEN "1001" => SEG7 <= "0010000";	-- 9
		WHEN OTHERS => SEG7 <= "0000110";	-- E for Error
		END CASE;
	END PROCESS;

END BEHAVIOURAL;

